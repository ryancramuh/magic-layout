magic
tech sky130A
timestamp 1759298223
<< locali >>
rect 0 25 20 45
rect 390 25 410 45
<< metal1 >>
rect 0 220 20 310
rect 0 65 20 155
use inverter  inverter_0
timestamp 1759297225
transform 1 0 125 0 1 60
box -125 -55 80 275
use inverter  inverter_1
timestamp 1759297225
transform 1 0 330 0 1 60
box -125 -55 80 275
<< end >>
