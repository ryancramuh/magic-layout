magic
tech sky130A
timestamp 1759800970
<< nwell >>
rect -120 135 85 390
<< nmos >>
rect 0 0 15 100
<< pmos >>
rect 0 155 15 370
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
<< pdiff >>
rect -50 355 0 370
rect -50 285 -35 355
rect -15 285 0 355
rect -50 240 0 285
rect -50 170 -35 240
rect -15 170 0 240
rect -50 155 0 170
rect 15 355 65 370
rect 15 285 30 355
rect 50 285 65 355
rect 15 240 65 285
rect 15 170 30 240
rect 50 170 65 240
rect 15 155 65 170
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
<< pdiffc >>
rect -35 285 -15 355
rect -35 170 -15 240
rect 30 285 50 355
rect 30 170 50 240
<< psubdiff >>
rect -100 85 -50 100
rect -100 15 -85 85
rect -65 15 -50 85
rect -100 0 -50 15
<< nsubdiff >>
rect -100 355 -50 370
rect -100 285 -85 355
rect -65 285 -50 355
rect -100 240 -50 285
rect -100 170 -85 240
rect -65 170 -50 240
rect -100 155 -50 170
<< psubdiffcont >>
rect -85 15 -65 85
<< nsubdiffcont >>
rect -85 285 -65 355
rect -85 170 -65 240
<< poly >>
rect 0 370 15 385
rect 0 140 15 155
rect 0 100 15 115
rect 0 -15 15 0
<< locali >>
rect -100 405 -70 410
rect -100 385 -95 405
rect -75 385 -70 405
rect -100 365 -70 385
rect -100 355 -5 365
rect -100 285 -85 355
rect -65 285 -35 355
rect -15 285 -5 355
rect -100 275 -5 285
rect 20 355 65 365
rect 20 285 30 355
rect 50 285 65 355
rect 20 275 65 285
rect -100 240 -5 250
rect -100 170 -85 240
rect -65 170 -35 240
rect -15 170 -5 240
rect -100 160 -5 170
rect 20 240 65 250
rect 20 170 30 240
rect 50 170 65 240
rect 20 160 65 170
rect -100 135 -75 160
rect -120 115 -75 135
rect 20 135 45 160
rect 20 115 85 135
rect 20 95 45 115
rect -100 85 -5 95
rect -100 15 -85 85
rect -65 15 -35 85
rect -15 15 -5 85
rect -100 5 -5 15
rect 20 85 65 95
rect 20 15 30 85
rect 50 15 65 85
rect 20 5 65 15
rect -100 -10 -70 5
rect -100 -30 -95 -10
rect -75 -30 -70 -10
rect -100 -40 -70 -30
<< viali >>
rect -95 385 -75 405
rect -95 -30 -75 -10
<< metal1 >>
rect -120 405 85 410
rect -120 385 -95 405
rect -75 385 85 405
rect -120 375 85 385
rect -120 -10 85 -5
rect -120 -30 -95 -10
rect -75 -30 85 -10
rect -120 -40 85 -30
<< labels >>
flabel locali -120 125 -120 125 3 FreeSans 320 0 0 0 A
port 1 e
flabel locali 85 125 85 125 7 FreeSans 320 0 0 0 Y
port 2 w
flabel metal1 85 395 85 395 7 FreeSans 320 0 0 0 VP
port 3 w
flabel metal1 85 -25 85 -25 7 FreeSans 320 0 0 0 VN
port 4 w
rlabel locali 65 215 65 215 3 B
<< end >>
